module ball(input logic clk,
	input logic reset_n,
	output logic );



endmodule // ball